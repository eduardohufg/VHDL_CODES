LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


ENTITY CONTACOMP IS
	PORT(CLK, RST, START: IN STD_LOGIC;
			S: OUT STD_LOGIC_VECTOR (4 DOWNTO 0));
			
	END CONTACOMP;
	
	
ARCHITECTURE RTL OF CONTACOMP IS

	COMPONENT CONTADOR24BITS IS
	PORT(CLK, RST, START: IN STD_LOGIC;
			O: OUT STD_LOGIC);
	END  COMPONENT CONTADOR24BITS;
	

	COMPONENT CONTADOR5BITS IS 
	PORT(ENA,CLK, RST: IN STD_LOGIC;
			S: OUT STD_LOGIC_VECTOR(4 DOWNTO 0));
	
	END COMPONENT CONTADOR5BITS;
	
	SIGNAL OV: STD_LOGIC;
	
	
	BEGIN
	
		I0: CONTADOR24BITS PORT MAP(CLK, RST, START, OV);
		
		I1: CONTADOR5BITS PORT MAP(OV, CLK, RST, S);
		
	END RTL;