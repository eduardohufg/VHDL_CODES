LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


ENTITY LCD IS
	PORT(CLK, RST, START: IN STD_LOGIC;
			E, RS, RW, LCD_BLON, LCD_ON: OUT STD_LOGIC;
			DATA: OUT STD_LOGIC_VECTOR (7 DOWNTO 0));
	END LCD;
	
	
ARCHITECTURE RTL OF LCD IS

	COMPONENT CONTADOR15BITS IS
		PORT(CLK, RST, START: IN STD_LOGIC; --Bits de control
				O: OUT STD_LOGIC); --Over Flow del contador
	END COMPONENT CONTADOR15BITS;
	
	COMPONENT MESTADOSLCD IS

	PORT (
		CLK, RST, ENA_LCD : IN STD_LOGIC;
		RS, RW, E, LCD_BLON, LCD_ON : OUT STD_LOGIC;
		DATA : OUT STD_LOGIC_VECTOR (7 DOWNTO 0));
	
	END COMPONENT MESTADOSLCD;
	
	
	SIGNAL OV: STD_LOGIC;
	
	BEGIN 
		
		IO: CONTADOR15BITS PORT MAP(CLK, RST,START, OV);
		I1: MESTADOSLCD PORT MAP (CLK, RST, OV, RS, RW, E, LCD_BLON, LCD_ON, DATA);
		
	END RTL;