LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY SUMA_MULT_4S IS
	PORT (COEF: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
				B_3: IN STD_LOGIC;
				M: OUT STD_LOGIC_VECTOR(8 DOWNTO 0));
	END SUMA_MULT_4S;
	
ARCHITECTURE RTL OF SUMA_MULT_4S IS
	COMPONENT ha IS

		PORT (a,b : IN STD_LOGIC;
      s, Cout: OUT STD_LOGIC);
	END COMPONENT ha;
	
	COMPONENT fa IS

		PORT (a,b, Cin : IN STD_LOGIC;
      s, Cout: OUT STD_LOGIC);
	END COMPONENT fa;

SIGNAL C: STD_LOGIC_VECTOR(15 DOWNTO 1);
SIGNAL S: STD_LOGIC_VECTOR(9 DOWNTO 1);

BEGIN

M(0) <= COEF(0);


I0: ha port map (COEF(1), COEF(4), M(1), C(1));
I1: FA PORT MAP (COEF(2), COEF(5), C(1), S(1), C(2));
I2: FA PORT MAP (COEF(3), COEF(6), C(2), S(2), C(3));
I3: FA PORT MAP (COEF(3), COEF(7), C(3), S(3), C(4));
I4: FA PORT MAP (COEF(3), COEF(7), C(4), S(4), C(5));
I5: FA PORT MAP (COEF(3), COEF(7), C(5), S(5), C(6));


I6: HA PORT MAP (COEF(8), S(1), M(2), C(7));
I7: FA PORT MAP (COEF(9), S(2), C(7), S(6), C(8));
I8: FA PORT MAP (COEF(10), S(3), C(8), S(7), C(9));
I9: FA PORT MAP (COEF(11), S(4), C(9), S(8), C(10));
I10: FA PORT MAP (COEF(11), S(5), C(10), S(9), C(11));


I11: FA PORT MAP(COEF(12), S(6), B_3, M(3), C(12));
I12: FA PORT MAP(COEF(13), S(7), C(12), M(4), C(13));
I13: FA PORT MAP(COEF(14), S(8), C(13), M(5), C(14));
I14: FA PORT MAP(COEF(15), S(9), C(14), M(6), C(15));

I15: FA PORT MAP(C(6), C(11), C(15), M(7), M(8));

END RTL;


 






