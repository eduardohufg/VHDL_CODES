--Circuio: Detector de secuencia de 4 bits--
--Autor: Eduardo Chavez Martin A01799595--


LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY DET_SEQ_4BITS IS
	PORT (CLK, RST, I: IN STD_LOGIC;
			ESTATOS: OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
			O: OUT STD_LOGIC);
			
	END DET_SEQ_4BITS;
	
ARCHITECTURE RTL OF DET_SEQ_4BITS IS
	TYPE EDOS IS (IDLE, E1 ,E2, E3, E4);
	
	SIGNAL EDO, EDOF : EDOS;
BEGIN

P1: PROCESS (CKL, RST) IS
	BEGIN
		IF(RST = '0') THEN
			EDO <= IDLE;
		ELSIF (CLK 'EVENT AND CLK = '1') THEN
			EDO <= EDOF;
		END IF
END PROCESS P1;

P2: PROCESS (EDO, I) IS
BEGIN 
	CASE EDO IS
		WHEN IDLE => IF(I = '0') THEN
							EDOF <= IDLE;
						ELSE 
							


	
