LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY SUMA_MULT4 IS
	PORT( A, B: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
			M: OUT STD_LOGIC_VECTOR(8 DOWNTO 0));
			
	END SUMA_MULT4;
	
ARCHITECTURE RTL OF SUMA_MULT4 IS

	
	COMPONENT CODER_4_S is
		Port ( A,B : in  STD_LOGIC_VECTOR (3 downto 0);
           COEF : out  STD_LOGIC_VECTOR (15 downto 0));
	end COMPONENT CODER_4_S;

	COMPONENT SUMA_MULT_4S IS
	PORT (COEF: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
				B_3: IN STD_LOGIC;
				M: OUT STD_LOGIC_VECTOR(8 DOWNTO 0));
	END COMPONENT SUMA_MULT_4S;

SIGNAL COEF: STD_LOGIC_VECTOR(15 DOWNTO 0);

BEGIN 

I0: CODER_4_S PORT MAP(A,B, COEF);
I1: SUMA_MULT_4S PORT MAP(COEF, B(3), M);

END RTL;
