--Circuito: Sumador BCD de dos digitos
--Autor: Eduardo Chavez Martin A01799595
-- Curso: TE2002B --

-- Seccion de definicion de Librerias --

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
--Declaramos entidad

ENTITY BCD_8BITS IS
	PORT (DATO: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
			S1,S2: IN STD_LOGIC;
			SALIDA: OUT STD_LOGIC_VECTOR(13 DOWNTO 0));
	END BCD_8BITS;
--Arquitecruta
	
ARCHITECTURE ARC OF BCD_8BITS IS
	
	--Descripcion de los componentes a utilizar
	COMPONENT SUM_BCD IS
	PORT(A,B: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
			CIN: IN STD_LOGIC;
			S: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
			COUT: OUT STD_LOGIC);
		END COMPONENT SUM_BCD;
	
	COMPONENT BIN2BCD IS
	PORT(BIN: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
			BCD: OUT STD_LOGIC_VECTOR (3 DOWNTO 0));
		END COMPONENT BIN2BCD;
		
	COMPONENT BCD_CODER IS
	PORT(BCD: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			SEG: OUT STD_LOGIC_VECTOR (6 DOWNTO 0));
		END COMPONENT BCD_CODER;
		
	--Signals para conectar y almacenar datos
	SIGNAL BC1: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL SIG1, SIG2: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL CO1, CO2: STD_LOGIC;
	SIGNAL SUM1, SUM2: STD_LOGIC_VECTOR (3 DOWNTO 0);
	SIGNAL SAL1: STD_LOGIC_VECTOR (13 DOWNTO 0);
	BEGIN
		
		I0: BIN2BCD PORT MAP(DATO(3 DOWNTO 0), BC1(3 DOWNTO 0));
		I1: BIN2BCD PORT MAP(DATO(7 DOWNTO 4), BC1(7 DOWNTO 4));
	
	--Procesos para la asignacion de datos a los registros
		PROCESS (S1)
			BEGIN
			
				IF S1 = '1' THEN 
					SIG1 <= BC1;
				END IF;
			END PROCESS;
			
		PROCESS (S2)
			BEGIN 
		
			IF S2 = '1' THEN
				SIG2 <= BC1;
			END IF;
		END PROCESS;
			
		--Mapeo y conexion de los componentes
		I2: SUM_BCD PORT MAP(SIG1(3 DOWNTO 0), SIG2(3 DOWNTO 0),'0', SUM1, CO1);
		I3: SUM_BCD PORT MAP(SIG1(7 DOWNTO 4), SIG2(7 DOWNTO 4), CO1, SUM2, CO2);
		
		I4: BCD_CODER PORT MAP(SUM1, SAL1(6 DOWNTO 0));
		I5: BCD_CODER PORT MAP(SUM2, SAL1(13 DOWNTO 7));
		
		SALIDA <= SAL1;
		END ARC;
		
			
			
			
			
			