LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;


ENTITY BIN2GR IS 
	PORT (INP: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
			SEL: IN STD_LOGIC;
			S: OUT STD_LOGIC_VECTOR(2 DOWNTO 0));
	END BIN2GR;
	
ARCHITECTURE ARC OF BIN2GR IS

BEGIN

	S(2) <= INP(2);
	S(1) <= INP(2) XOR INP(1);
	
	S(0) <= (INP(1) XOR INP(0)) WHEN SEL = '0' ELSE
				(INP(2) XOR INP(1) XOR INP(0));

END ARC;