--Circuio: Generador de secuencia de 3 bits--
--Autor: Eduardo Chavez Martin A01799595--
--Curso: TE2002B

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY SECUENCIA_3BITS IS 
PORT (CLK, RST: IN STD_LOGIC;
		SALIDA: OUT STD_LOGIC_VECTOR (2 DOWNTO 0));
		END SECUENCIA_3BITS;
		
ARCHITECTURE RTL OF SECUENCIA_3BITS IS

SIGNAL EDO,EDOF: STD_LOGIC_VECTOR(2 DOWNTO 0);

BEGIN 

P1: PROCESS (CLK,RST) IS

BEGIN 
	IF(RST = '0') THEN
		EDO<="000";
	ELSIF (CLK'EVENT AND CLK = '1') THEN
		EDO <= EDOF;
	END IF;
END PROCESS P1;


--DEFINIR LAS TRANCISIONES DEL AUTOMATA

P2: PROCESS (EDO)
	BEGIN
	
		CASE EDO IS
			WHEN "000" => EDOF <= "100";
			WHEN "010" => EDOF <= "011";
			WHEN "011" => EDOF <= "000";
			WHEN "100" => EDOF <= "111";
			WHEN "111" => EDOF <= "010";
			WHEN OTHERS => NULL;
		END CASE;
	END PROCESS P2;
	
	SALIDA <= EDO;  --CONECTANDO LAS SALIDAS A LOS FLIPFLOPS D
	
END RTL;

